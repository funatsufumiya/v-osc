// Package osc provides a package for sending and receiving OpenSoundControl
// messages. The package is implemented in pure Go.
module osc

import net
import time

// import (
// 	"bufio"
// 	"bytes"
// 	"encoding"
// 	"encoding/binary"
// 	"errors"
// 	"fmt"
// 	"net"
// 	"reflect"
// 	"regexp"
// 	"strings"
// 	"time"
// )

const secondsFrom1900To1970  = 2208988800                      // Source: RFC 868
const nanosecondsPerFraction = f64(0.23283064365386962891)    // 1e9/(2^32)
const bundleTagString       = "#bundle"

// Packet is the interface for Message and Bundle.
pub interface Packet {
	encoding.BinaryMarshaler
}

// Message represents a single OSC message. An OSC message consists of an OSC
// address pattern and zero or more arguments.
pub struct Message {
pub mut:
	address   string
	arguments []interface{}
}

// Verify that Messages implements the Packet interface.
var _ Packet = (*Message)(nil)

// Bundle represents an OSC bundle. It consists of the OSC-string "#bundle"
// followed by an OSC Time Tag, followed by zero or more OSC bundle/message
// elements. The OSC-timetag is a 64-bit fixed point time tag. See
// http://opensoundcontrol.org/spec-1_0 for more information.
pub struct Bundle {
pub mut:
	timetag  Timetag
	messages []*Message
	bundles  []*Bundle
}

// Verify that Bundle implements the Packet interface.
var _ Packet = (*Bundle)(nil)

// Client enables you to send OSC packets. It sends OSC messages and bundles to
// the given IP address and port.
pub struct Client {
	ip    string
	port  int
	laddr *net.UDPAddr
}

// Server represents an OSC server. The server listens on Address and Port for
// incoming OSC packets and bundles.
pub struct Server {
pub mut:
	addr        string
	dispatcher  Dispatcher
	read_timeout time.Duration
	close       func() error
}

// Timetag represents an OSC Time Tag.
// An OSC Time Tag is defined as follows:
// Time tags are represented by a 64 bit fixed point number. The first 32 bits
// specify the number of seconds since midnight on January 1, 1900, and the
// last 32 bits specify fractional parts of a second to a precision of about
// 200 picoseconds. This is the representation used by Internet NTP timestamps.
pub struct Timetag {
pub mut:
	time_tag  uint64 // The acutal time tag
	time     time.Time
	min_value uint64 // Minimum value of an OSC Time Tag. Is always 1.
}

// Dispatcher is an interface for an OSC message dispatcher. A dispatcher is
// responsible for dispatching received OSC messages.
interface Dispatcher {
	Dispatch(packet Packet)
}

// Handler is an interface for message handlers. Every handler implementation
// for an OSC message must implement this interface.
interface Handler {
	HandleMessage(msg *Message)
}

// HandlerFunc implements the Handler interface. Type definition for an OSC
// handler function.
type HandlerFunc func(msg *Message)

// HandleMessage calls itself with the given OSC Message. Implements the
// Handler interface.
fn (f HandlerFunc) handle_message(msg *Message) {
	f(msg)
}

////
// StandardDispatcher
////

// StandardDispatcher is a dispatcher for OSC packets. It handles the dispatching of
// received OSC packets to Handlers for their given address.
pub struct StandardDispatcher {
	handlers       map[string]Handler
	defaultHandler Handler
}

// NewStandardDispatcher returns an StandardDispatcher.
pub fn new_standard_dispatcher() *StandardDispatcher {
	return &StandardDispatcher{handlers: make(map[string]Handler)}
}

// AddMsgHandler adds a new message handler for the given OSC address.
pub fn (s *StandardDispatcher) add_msg_handler(addr string, handler HandlerFunc) error {
	if addr == "*" {
		s.defaultHandler = handler
		return nil
	}
	for _, chr := range "*?,[]{}# " {
		if strings.Contains(addr, fmt.Sprintf("%c", chr)) {
			return errors.new("OSC Address string may not contain any characters in \"*?,[]{}#")
		}
	}

	if address_exists(addr, s.handlers) {
		return errors.new("OSC address exists already")
	}

	s.handlers[addr] = handler
	return nil
}

// Dispatch dispatches OSC packets. Implements the Dispatcher interface.
pub fn (s *StandardDispatcher) dispatch(packet Packet) {
	switch p := packet.(type) {
	default:
		return

	case *Message:
		for addr, handler := range s.handlers {
			if p.matches(addr) {
				handler.handle_message(p)
			}
		}
		if s.defaultHandler != nil {
			s.defaultHandler.handle_message(p)
		}

	case *Bundle:
		timer := time.new_timer(p.Timetag.expires_in())

		go func() {
			<-timer.C
			for _, message := range p.Messages {
				for address, handler := range s.handlers {
					if message.matches(address) {
						handler.handle_message(message)
					}
				}
				if s.defaultHandler != nil {
					s.defaultHandler.handle_message(message)
				}
			}

			// Process all bundles
			for _, b := range p.Bundles {
				s.dispatch(b)
			}
		}()
	}
}

////
// Message
////

// NewMessage returns a new Message. The address parameter is the OSC address.
pub fn new_message(addr string, args ...interface{}) *Message {
	return &Message{Address: addr, Arguments: args}
}

// Append appends the given arguments to the arguments list.
pub fn (msg *Message) append(args ...interface{}) {
	msg.Arguments = append(msg.Arguments, args...)
}

// Equals returns true if the given OSC Message `m` is equal to the current OSC
// Message. It checks if the OSC address and the arguments are equal. Returns
// true if the current object and `m` are equal.
pub fn (msg *Message) equals(m *Message) bool {
	return reflect.deep_equal(msg, m)
}

// Clear clears the OSC address and all arguments.
pub fn (msg *Message) clear() {
	msg.Address = ""
	msg.ClearData()
}

// ClearData removes all arguments from the OSC Message.
pub fn (msg *Message) clear_data() {
	msg.Arguments = msg.arguments[len(msg.Arguments):]
}

// matches returns true, if the OSC address pattern of the OSC Message matches the given
// address. The match is case sensitive!
pub fn (msg *Message) matches(addr string) bool {
	exp := get_reg_ex(msg.Address)
	return exp.matches_string(addr)
}

// TypeTags returns the type tag string.
pub fn (msg *Message) type_tags() (string, error) {
	if msg == nil {
		return "", fmt.Errorf("message is nil")
	}

	tags := ","
	for _, m := range msg.Arguments {
		s, err := get_type_tag(m)
		if err != nil {
			return "", err
		}
		tags += s
	}

	return tags, nil
}

// String implements the fmt.Stringer interface.
pub fn (msg *Message) String() string {
	if msg == nil {
		return ""
	}

	tags, err := msg.type_tags()
	if err != nil {
		return ""
	}

	formatString := "%s %s"
	var args []interface{}
	args = append(args, msg.Address)
	args = append(args, tags)

	for _, arg := range msg.Arguments {
		switch arg.(type) {
		case bool, int32, int64, float32, float64, string:
			formatString += " %v"
			args = append(args, arg)

		case nil:
			formatString += " %s"
			args = append(args, "Nil")

		case []byte:
			formatString += " %s"
			args = append(args, "blob")

		case Timetag:
			formatString += " %d"
			timeTag := arg.(Timetag)
			args = append(args, timeTag.time_tag())
		}
	}

	return fmt.Sprintf(formatString, args...)
}

// CountArguments returns the number of arguments.
pub fn (msg *Message) count_arguments() int {
	return len(msg.Arguments)
}

// MarshalBinary serializes the OSC message to a byte buffer. The byte buffer
// has the following format:
// 1. OSC Address Pattern
// 2. OSC Type Tag String
// 3. OSC Arguments
pub fn (msg *Message) marshal_binary() ([]byte, error) {
	// We can start with the OSC address and add it to the buffer
	data := new(bytes.Buffer)
	if _, err := write_padded_string(msg.Address, data); err != nil {
		return nil, err
	}

	// Type tag string starts with ","
	typetags := []byte{','}

	// Process the type tags and collect all arguments
	payload := new(bytes.Buffer)
	for _, arg := range msg.Arguments {
		// FIXME: Use t instead of arg
		switch t := arg.(type) {
		default:
			return nil, fmt.Errorf("OSC - unsupported type: %T", t)

		case bool:
			if arg.(bool) {
				typetags = append(typetags, 'T')
			} else {
				typetags = append(typetags, 'F')
			}

		case nil:
			typetags = append(typetags, 'N')

		case int32:
			typetags = append(typetags, 'i')
			if err := binary.write(payload, binary.BigEndian, int32(t)); err != nil {
				return nil, err
			}

		case float32:
			typetags = append(typetags, 'f')
			if err := binary.write(payload, binary.BigEndian, float32(t)); err != nil {
				return nil, err
			}

		case string:
			typetags = append(typetags, 's')
			if _, err := write_padded_string(t, payload); err != nil {
				return nil, err
			}

		case []byte:
			typetags = append(typetags, 'b')
			if _, err := write_blob(t, payload); err != nil {
				return nil, err
			}

		case int64:
			typetags = append(typetags, 'h')
			if err := binary.write(payload, binary.BigEndian, int64(t)); err != nil {
				return nil, err
			}

		case float64:
			typetags = append(typetags, 'd')
			if err := binary.write(payload, binary.BigEndian, float64(t)); err != nil {
				return nil, err
			}

		case Timetag:
			typetags = append(typetags, 't')
			timeTag := arg.(Timetag)
			b, err := timeTag.marshal_binary()
			if err != nil {
				return nil, err
			}
			if _, err = payload.write(b); err != nil {
				return nil, err
			}
		}
	}

	// Write the type tag string to the data buffer
	if _, err := write_padded_string(string(typetags), data); err != nil {
		return nil, err
	}

	// Write the payload (OSC arguments) to the data buffer
	if _, err := data.write(payload.bytes()); err != nil {
		return nil, err
	}

	return data.bytes(), nil
}

////
// Bundle
////

// NewBundle returns an OSC Bundle. Use this function to create a new OSC
// Bundle.
pub fn new_bundle(time time.Time) *Bundle {
	return &Bundle{Timetag: *new_timetag(time)}
}

// Append appends an OSC bundle or OSC message to the bundle.
pub fn (b *Bundle) append(pck Packet) error {
	switch t := pck.(type) {
	default:
		return fmt.Errorf("unsupported OSC packet type: only Bundle and Message are supported")

	case *Bundle:
		b.Bundles = append(b.Bundles, t)

	case *Message:
		b.Messages = append(b.Messages, t)
	}

	return nil
}

// MarshalBinary serializes the OSC bundle to a byte array with the following
// format:
// 1. Bundle string: '#bundle'
// 2. OSC timetag
// 3. Length of first OSC bundle element
// 4. First bundle element
// 5. Length of n OSC bundle element
// 6. n bundle element
pub fn (b *Bundle) marshal_binary() ([]byte, error) {
	// Add the '#bundle' string
	data := new(bytes.Buffer)
	if _, err := write_padded_string("#bundle", data); err != nil {
		return nil, err
	}

	// Add the time tag
	bd, err := b.Timetag.marshal_binary()
	if err != nil {
		return nil, err
	}
	if _, err = data.write(bd); err != nil {
		return nil, err
	}

	// Process all OSC Messages
	for _, m := range b.Messages {
		buf, err := m.marshal_binary()
		if err != nil {
			return nil, err
		}

		// Append the length of the OSC message
		if err = binary.write(data, binary.BigEndian, int32(len(buf))); err != nil {
			return nil, err
		}

		// Append the OSC message
		if _, err = data.write(buf); err != nil {
			return nil, err
		}
	}

	// Process all OSC Bundles
	for _, b := range b.Bundles {
		buf, err := b.marshal_binary()
		if err != nil {
			return nil, err
		}

		// Write the size of the bundle
		if err = binary.write(data, binary.BigEndian, int32(len(buf))); err != nil {
			return nil, err
		}

		// Append the bundle
		_, err = data.write(buf)
		if err != nil {
			return nil, err
		}
	}

	return data.bytes(), nil
}

////
// Client
////

// NewClient creates a new OSC client. The Client is used to send OSC
// messages and OSC bundles over an UDP network connection. The `ip` argument
// specifies the IP address and `port` defines the target port where the
// messages and bundles will be send to.
pub fn new_client(ip string, port int) *Client {
	return &Client{ip: ip, port: port, laddr: nil}
}

// IP returns the IP address.
pub fn (c *Client) ip() string { return c.ip }

// SetIP sets a new IP address.
pub fn (c *Client) set_ip(ip string) { c.ip = ip }

// Port returns the port.
pub fn (c *Client) port() int { return c.port }

// SetPort sets a new port.
pub fn (c *Client) set_port(port int) { c.port = port }

// SetLocalAddr sets the local address.
pub fn (c *Client) set_local_addr(ip string, port int) error {
	laddr, err := net.resolve_udpaddr("udp", fmt.Sprintf("%s:%d", ip, port))
	if err != nil {
		return err
	}
	c.laddr = laddr
	return nil
}

// Send sends an OSC Bundle or an OSC Message.
pub fn (c *Client) send(packet Packet) error {
	addr, err := net.resolve_udpaddr("udp", fmt.Sprintf("%s:%d", c.ip, c.port))
	if err != nil {
		return err
	}
	conn, err := net.dial_udp("udp", c.laddr, addr)
	if err != nil {
		return err
	}
	defer conn.close()

	data, err := packet.marshal_binary()
	if err != nil {
		return err
	}

	if _, err = conn.write(data); err != nil {
		return err
	}
	return nil
}

////
// Server
////

// ListenAndServe retrieves incoming OSC packets and dispatches the retrieved
// OSC packets.
pub fn (s *Server) listen_and_serve() error {
	defer s.close_connection()

	if s.Dispatcher == nil {
		s.Dispatcher = new_standard_dispatcher()
	}

	ln, err := net.listen_packet("udp", s.Addr)
	if err != nil {
		return err
	}

	s.close = ln.Close

	return s.serve(ln)
}

// Serve retrieves incoming OSC packets from the given connection and dispatches
// retrieved OSC packets. If something goes wrong an error is returned.
pub fn (s *Server) serve(c net.PacketConn) error {
	var tempDelay time.Duration
	for {
		msg, err := s.read_from_connection(c)
		if err != nil {
			if ne, ok := err.(net.error); ok && ne.temporary() {
				if tempDelay == 0 {
					tempDelay = 5 * time.millisecond
				} else {
					tempDelay *= 2
				}
				if max := 1 * time.second; tempDelay > max {
					tempDelay = max
				}
				time.Sleep(tempDelay)
				continue
			}
			return err
		}
		tempDelay = 0
		go s.Dispatcher.dispatch(msg)
	}
}

// CloseConnection forcibly closes a server's connection.
//
// This causes a "use of closed network connection" error the next time the
// server attempts to read from the connection.
pub fn (s *Server) close_connection() error {
	if s.close == nil {
		return nil
	}

	err := s.close()
	// If we get "use of closed network connection", it's not a problem because
	// closing the network connection is exactly what we wanted to do!
	if err != nil && !strings.contains(
		err.Error(), "use of closed network connection",
	) {
		return err
	}

	return nil
}

// ReceivePacket listens for incoming OSC packets and returns the packet if one is received.
pub fn (s *Server) receive_packet(c net.PacketConn) (Packet, error) {
	return s.read_from_connection(c)
}

// readFromConnection retrieves OSC packets.
fn (s *Server) read_from_connection(c net.PacketConn) (Packet, error) {
	if s.ReadTimeout != 0 {
		if err := c.set_read_deadline(time.now().add(s.read_timeout)); err != nil {
			return nil, err
		}
	}

	data := make([]byte, 65535)
	n, _, err := c.read_from(data)
	if err != nil {
		return nil, err
	}

	p, err := read_packet(bufio.new_reader(bytes.new_buffer(data[0:n])))
	if err != nil {
		return nil, err
	}
	return p, nil
}

// ParsePacket parses the given msg string and returns a Packet
pub fn parse_packet(msg string) (Packet, error) {
	p, err := read_packet(bufio.new_reader(bytes.new_bufferString(msg)))
	if err != nil {
		return nil, err
	}
	return p, nil
}

// receivePacket receives an OSC packet from the given reader.
fn read_packet(reader *bufio.Reader) (Packet, error) {
	//var buf []byte
	buf, err := reader.Peek(1)
	if err != nil {
		return nil, err
	}

	// An OSC Message starts with a '/'
	if buf[0] == '/' {
		packet, err := read_message(reader)
		if err != nil {
			return nil, err
		}
		return packet, nil
	}
	if buf[0] == '#' { // An OSC bundle starts with a '#'
		packet, err := read_bundle(reader)
		if err != nil {
			return nil, err
		}
		return packet, nil
	}

	var p Packet
	return p, nil
}

// readBundle reads an Bundle from reader.
fn read_bundle(reader *bufio.Reader) (*Bundle, error) {
	// Read the '#bundle' OSC string
	startTag, _, err := read_padded_string(reader)
	if err != nil {
		return nil, err
	}

	if startTag != bundle_tag_string {
		return nil, fmt.Errorf("invalid bundle start tag: %s", startTag)
	}

	// Read the timetag
	var timeTag uint64
	if err := binary.read(reader, binary.big_endian, &timeTag); err != nil {
		return nil, err
	}

	// Create a new bundle
	bundle := new_bundle(timetag_to_time(timeTag))

	// Read until the end of the buffer
	for reader.buffered() > 0 {
		// Read the size of the bundle element
		var length int32
		if err := binary.read(reader, binary.big_endian, &length); err != nil {
			return nil, err
		}

		p, err := read_packet(reader)
		if err != nil {
			return nil, err
		}
		if err = bundle.append(p); err != nil {
			return nil, err
		}
	}

	return bundle, nil
}

// readMessage from `reader`.
fn read_message(reader *bufio.Reader) (*Message, error) {
	// First, read the OSC address
	addr, _, err := read_padded_string(reader)
	if err != nil {
		return nil, err
	}

	// Read all arguments
	msg := new_message(addr)
	if err = read_arguments(msg, reader); err != nil {
		return nil, err
	}

	return msg, nil
}

// readArguments from `reader` and add them to the OSC message `msg`.
fn read_arguments(msg *Message, reader *bufio.Reader) error {
	// Read the type tag string
	typetags, _, err := read_padded_string(reader)
	if err != nil {
		return err
	}

	if len(typetags) == 0 {
		return nil
	}

	// If the typetag doesn't start with ',', it's not valid
	if typetags[0] != ',' {
		return fmt.Errorf("unsupported type tag string %s", typetags)
	}

	// Remove ',' from the type tag
	typetags = typetags[1:]

	for _, c := range typetags {
		switch c {
		default:
			return fmt.Errorf("unsupported type tag: %c", c)

		case 'i': // int32
			var i int32
			if err = binary.read(reader, binary.BigEndian, &i); err != nil {
				return err
			}
			msg.append(i)

		case 'h': // int64
			var i int64
			if err = binary.read(reader, binary.BigEndian, &i); err != nil {
				return err
			}
			msg.append(i)

		case 'f': // float32
			var f float32
			if err = binary.read(reader, binary.BigEndian, &f); err != nil {
				return err
			}
			msg.append(f)

		case 'd': // float64/double
			var d float64
			if err = binary.read(reader, binary.BigEndian, &d); err != nil {
				return err
			}
			msg.append(d)

		case 's': // string
			// TODO: fix reading string value
			var s string
			if s, _, err = read_padded_string(reader); err != nil {
				return err
			}
			msg.append(s)

		case 'b': // blob
			var buf []byte
			if buf, _, err = read_blob(reader); err != nil {
				return err
			}
			msg.append(buf)

		case 't': // OSC time tag
			var tt uint64
			if err = binary.read(reader, binary.big_endian, &tt); err != nil {
				return nil
			}
			msg.append(*new_timetag_from_timetag(tt))

		case 'N': // nil
			msg.append(nil)

		case 'T': // true
			msg.append(true)

		case 'F': // false
			msg.append(false)
		}
	}

	return nil
}

////
// Timetag
////

// NewTimetag returns a new OSC time tag object.
pub fn new_timetag(ts time.Time) *Timetag {
	return &Timetag{
		time:     ts,
		timeTag:  time_to_timetag(ts),
		MinValue: uint64(1)}
}

// NewTimetagFromTimetag creates a new Timetag from the given `timetag`.
pub fn new_timetag_from_timetag(timetag uint64) *Timetag {
	time := timetag_to_time(timetag)
	return new_timetag(time)
}

// Time returns the time.
pub fn (t *Timetag) time() time.Time {
	return t.time
}

// FractionalSecond returns the last 32 bits of the OSC time tag. Specifies the
// fractional part of a second.
pub fn (t *Timetag) fractional_second() uint32 {
	return uint32(t.timeTag << 32)
}

// SecondsSinceEpoch returns the first 32 bits (the number of seconds since the
// midnight 1900) from the OSC time tag.
pub fn (t *Timetag) seconds_since_epoch() uint32 {
	return uint32(t.timeTag >> 32)
}

// TimeTag returns the time tag value
pub fn (t *Timetag) time_tag() uint64 {
	return t.timeTag
}

// MarshalBinary converts the OSC time tag to a byte array.
pub fn (t *Timetag) marshal_binary() ([]byte, error) {
	data := new(bytes.Buffer)
	if err := binary.write(data, binary.big_endian, t.timeTag); err != nil {
		return []byte{}, err
	}
	return data.bytes(), nil
}

// SetTime sets the value of the OSC time tag.
pub fn (t *Timetag) set_time(time time.Time) {
	t.time = time
	t.timeTag = time_to_timetag(time)
}

// ExpiresIn calculates the number of seconds until the current time is the
// same as the value of the time tag. It returns zero if the value of the
// time tag is in the past.
pub fn (t *Timetag) expires_in() time.Duration {
	// If the timetag is one the OSC method must be invoke immediately.
	// See https://ccrma.stanford.edu/groups/osc/spec-1_0.html#timetags.
	if t.timeTag <= 1 {
		return 0
	}

	tt := timetag_to_time(t.timeTag)
	seconds := time.Until(tt)

	// Invoke the OSC method immediately if the timetag is before or equal to the current time
	if seconds <= 0 {
		return 0
	}

	return seconds
}

// timeToTimetag converts the given time to an OSC time tag.
//
// An OSC time tag is defined as follows:
// Time tags are represented by a 64 bit fixed point number. The first 32 bits
// specify the number of seconds since midnight on January 1, 1900, and the
// last 32 bits specify fractional parts of a second to a precision of about
// 200 picoseconds. This is the representation used by Internet NTP timestamps.
//
// The time tag value consisting of 63 zero bits followed by a one in the least
// significant bit is a special case meaning "immediately."
//
// See also https://ccrma.stanford.edu/groups/osc/spec-1_0.html#timetags.
fn time_to_timetag(v time.Time) (timetag uint64) {
	if v.is_zero() {
		// Means "immediately". It cannot occur otherwise as timetag == 0 gets
		// converted to January 1, 1900 while time.Time{} means year 1 in Go.
		// Use the IsZero method to detect it.
		return 1
	}

	seconds := uint64(v.Unix() + secondsFrom1900To1970)
	secondFraction := float64(v.nanosecond()) / nanosecondsPerFraction

	return (seconds << 32) + uint64(uint32(secondFraction))
}

// timetagToTime converts the given OSC timetag to a time object.
fn timetag_to_time(timetag uint64) (t time.Time) {
	// Special case when timetag is == 1 that means "immediately". In this case we return
	// the zero time instant.
	if timetag == 1 {
		return time.Time{}
	}

	seconds := int64(timetag>>32) - secondsFrom1900To1970
	nanoseconds := int64(nanosecondsPerFraction * float64(float64(timetag&(1<<32-1))))

	return time.Unix(
		seconds,
		nanoseconds,
	)
}

////
// De/Encoding functions
////

// readBlob reads an OSC blob from the blob byte array. Padding bytes are
// removed from the reader and not returned.
fn read_blob(reader *bufio.Reader) ([]byte, int, error) {
	// First, get the length
	var blobLen int32
	if err := binary.read(reader, binary.BigEndian, &blobLen); err != nil {
		return nil, 0, err
	}
	n := 4 + int(blobLen)

	if blobLen < 1 || blobLen > int32(reader.Buffered()) {
		return nil, 0, fmt.Errorf("readBlob: invalid blob length %d", blobLen)
	}

	// Read the data
	blob := make([]byte, blobLen)
	if _, err := reader.read(blob); err != nil {
		return nil, 0, err
	}

	// Remove the padding bytes
	numPadBytes := pad_bytes_needed(int(blobLen))
	if numPadBytes > 0 {
		n += numPadBytes
		dummy := make([]byte, numPadBytes)
		if _, err := reader.read(dummy); err != nil {
			return nil, 0, err
		}
	}

	return blob, n, nil
}

// writeBlob writes the data byte array as an OSC blob into buff. If the length
// of data isn't 32-bit aligned, padding bytes will be added.
fn write_blob(data []byte, buf *bytes.Buffer) (int, error) {
	// Add the size of the blob
	dlen := int32(len(data))
	if err := binary.write(buf, binary.BigEndian, dlen); err != nil {
		return 0, err
	}

	// Write the data
	if _, err := buf.write(data); err != nil {
		return 0, nil
	}

	// Add padding bytes if necessary
	numPadBytes := pad_bytes_needed(len(data))
	if numPadBytes > 0 {
		padBytes := make([]byte, numPadBytes)
		n, err := buf.write(padBytes)
		if err != nil {
			return 0, err
		}
		numPadBytes = n
	}

	return 4 + len(data) + numPadBytes, nil
}

// readPaddedString reads a padded string from the given reader. The padding
// bytes are removed from the reader.
fn read_padded_string(reader *bufio.Reader) (string, int, error) {
	// Read the string from the reader
	str, err := reader.read_string(0)
	if err != nil {
		return "", 0, err
	}
	n := len(str)

	// Remove the padding bytes (leaving the null delimiter)
	padLen := pad_bytes_needed(len(str))
	if padLen > 0 {
		n += padLen
		padBytes := make([]byte, padLen)
		if _, err = reader.read(padBytes); err != nil {
			return "", 0, err
		}
	}

	// Strip off the string delimiter
	return str[:len(str)-1], n, nil
}

// writePaddedString writes a string with padding bytes to the a buffer.
// Returns, the number of written bytes and an error if any.
fn write_padded_string(str string, buf *bytes.Buffer) (int, error) {
	// Truncate at the first null, just in case there is more than one present
	nullIndex := strings.Index(str, "\x00")
	if nullIndex > 0 {
		str = str[:nullIndex]
	}
	// Write the string to the buffer
	n, err := buf.write_string(str)
	if err != nil {
		return 0, err
	}

	// Always write a null terminator, as we stripped it earlier if it existed
	buf.write_byte(0)
	n++

	// Calculate the padding bytes needed and create a buffer for the padding bytes
	numPadBytes := pad_bytes_needed(n)
	if numPadBytes > 0 {
		padBytes := make([]byte, numPadBytes)
		// Add the padding bytes to the buffer
		n, err := buf.write(padBytes)
		if err != nil {
			return 0, err
		}
		numPadBytes = n
	}

	return n + numPadBytes, nil
}

// padBytesNeeded determines how many bytes are needed to fill up to the next 4
// byte length.
fn pad_bytes_needed(elementLen int) int {
	return ((4 - (elementLen % 4)) % 4)
}

////
// Utility and helper functions
////

// PrintMessage pretty prints an OSC message to the standard output.
pub fn print_message(msg *Message) {
	fmt.Println(msg)
}

// addressExists returns true if the OSC address `addr` is found in `handlers`.
fn address_exists(addr string, handlers map[string]Handler) bool {
	for h := range handlers {
		if h == addr {
			return true
		}
	}
	return false
}

// getRegEx compiles and returns a regular expression object for the given
// address `pattern`.
fn get_reg_ex(pattern string) *regexp.Regexp {
	for _, trs := range []struct {
		old, new string
	}{
		{".", `\.`}, // Escape all '.' in the pattern
		{"(", `\(`}, // Escape all '(' in the pattern
		{")", `\)`}, // Escape all ')' in the pattern
		{"*", ".*"}, // Replace a '*' with '.*' that matches zero or more chars
		{"{", "("},  // Change a '{' to '('
		{",", "|"},  // Change a ',' to '|'
		{"}", ")"},  // Change a '}' to ')'
		{"?", "."},  // Change a '?' to '.'
	} {
		pattern = strings.replace(pattern, trs.old, trs.new, -1)
	}

	return regexp.must_compile(pattern)
}

// getTypeTag returns the OSC type tag for the given argument.
fn get_type_tag(arg interface{}) (string, error) {
	switch t := arg.(type) {
	case bool:
		if arg.(bool) {
			return "T", nil
		}
		return "F", nil
	case nil:
		return "N", nil
	case int32:
		return "i", nil
	case float32:
		return "f", nil
	case string:
		return "s", nil
	case []byte:
		return "b", nil
	case int64:
		return "h", nil
	case float64:
		return "d", nil
	case Timetag:
		return "t", nil
	default:
		return "", fmt.Errorf("unsupported type: %T", t)
	}
}
