module osc

// import (
// 	"bufio"
// 	"bytes"
// 	"io"
// 	"math/rand"
// 	"net"
// 	"reflect"
// 	"strconv"
// 	"strings"
// 	"sync"
// 	"testing"
// 	"time"
// )

fn message_append_test() {
	oscAddress := "/address"
	message := new_message(oscAddress)
	assert message.Address == oscAddress

	message.append("string argument")
	message.append(123456789)
	message.append(true)

	assert message.CountArguments() == 3
}

fn message_equals_test() {
	msg1 := new_message("/address")
	msg2 := new_message("/address")
	msg1.append(1234)
	msg2.append(1234)
	msg1.append("test string")
	msg2.append("test string")

	assert msg1.equals(msg2)
}

fn message_typetags_test() {

	struct TestData {
		desc string
		msg  &Message
		tags string
		ok   bool
	}

	test_data := [
		TestData{"addr_only", new_message("/"), ",", true},
		TestData{"nil", new_message("/", nil), ",N", true},
		TestData{"bool_true", new_message("/", true), ",T", true},
		TestData{"bool_false", new_message("/", false), ",F", true},
		TestData{"int32", new_message("/", int32(1)), ",i", true},
		TestData{"int64", new_message("/", int64(2)), ",h", true},
		TestData{"float32", new_message("/", float32(3.0)), ",f", true},
		TestData{"float64", new_message("/", float64(4.0)), ",d", true},
		TestData{"string", new_message("/", "5"), ",s", true},
		TestData{"[]byte", new_message("/", `6`), ",b", true},
		TestData{"two_args", new_message("/", "123", int32(456)), ",si", true},
		TestData{"invalid_msg", nil, "", false},
		TestData{"invalid_arg", new_message("/foo/bar", 789), "", false},
	]

	for tt in test_data  {
		tags, err := tt.msg.TypeTags()
		if err != nil && tt.ok {
			assert false, "${tt.desc}: TypeTags() unexpected error: ${err}"
			continue
		}
		if err == nil && !tt.ok {
			assert false, "${tt.desc}: TypeTags() expected an error"
			continue
		}
		if !tt.ok {
			continue
		}
		if got, want := tags, tt.tags; got != want {
			assert false, "${tt.desc}: TypeTags() = '${got}', want = '${want}'"
		}
	}
}

fn message_string_test() {
	for _, tt := range []struct {
		desc string
		msg  *Message
		str  string
	}{
		{"nil", nil, ""},
		{"addr_only", new_message("/foo/bar"), "/foo/bar ,"},
		{"one_addr", new_message("/foo/bar", "123"), "/foo/bar ,s 123"},
		{"two_args", new_message("/foo/bar", "123", int32(456)), "/foo/bar ,si 123 456"},
	} {
		if got, want := tt.msg.String(), tt.str; got != want {
			assert false, "${tt.desc}: String() = '${got}', want = '${want}'"
		}
	}
}

fn add_msg_handler_test() {
	d := NewStandardDispatcher()
	err := d.AddMsgHandler("/address/test", func(msg *Message) {})
	if err != nil {
		assert false, "Expected that OSC address '/address/test' is valid"
	}
}

fn add_msg_handler_with_invalid_address_test() {
	d := NewStandardDispatcher()
	err := d.AddMsgHandler("/address*/test", func(msg *Message) {})
	if err == nil {
		assert false, "Expected error with '/address*/test'"
	}
}

// These tests stop the server by forcibly closing the connection, which causes
// a "use of closed network connection" error the next time we try to read from
// the connection. As a workaround, this wraps server.ListenAndServe() in an
// error-handling layer that doesn't consider "use of closed network connection"
// an error.
//
// Open question: is this desired behavior, or should server.serve return
// successfully in cases where it would otherwise throw this error?
fn serve_until_interrupted(server *Server) error {
	if err := server.ListenAndServe(); err != nil &&
		!strings.Contains(err.Error(), "use of closed network connection") {
		return err
	}

	return nil
}

fn server_message_dispatching_test(stringArgument string) {
	finish := make(chan bool)
	start := make(chan bool)
	done := sync.WaitGroup{}
	done.Add(2)

	port := 6677
	addr := "localhost:" + strconv.Itoa(port)

	d := NewStandardDispatcher()
	server := &Server{Addr: addr, Dispatcher: d}

	defer func() {
		if err := server.CloseConnection(); err != nil {
			t.Error(err)
		}
	}()

	if err := d.AddMsgHandler(
		"/address/test",
		func(msg *Message) {
			defer func() {
				server.CloseConnection()
				finish <- true
			}()

			if len(msg.Arguments) != 2 {
				t.Errorf("Argument length should be 2 and is: %d", len(msg.Arguments))
			}

			if msg.Arguments[0].(int32) != 1122 {
				t.Error("Argument should be 1122 and is: " + string(msg.Arguments[0].(int32)))
			}

			receivedString := msg.Arguments[1].(string)

			if len(receivedString) != len(stringArgument) {
				t.Errorf(
					"String argument length should be %d and is %d",
					len(stringArgument),
					len(receivedString),
				)
			} else if receivedString != stringArgument {
				t.Errorf(
					"Argument should be %s and is: %s", stringArgument, receivedString,
				)
			}
		},
	); err != nil {
		t.Error("Error adding message handler")
	}

	// Server goroutine
	go func() {
		start <- true

		if err := serveUntilInterrupted(server); err != nil {
			t.Errorf("error during Serve: %s", err.Error())
		}
	}()

	// Client goroutine
	go func() {
		timeout := time.After(5 * time.Second)
		select {
		case <-timeout:
		case <-start:
			time.Sleep(500 * time.Millisecond)
			client := NewClient("localhost", port)
			msg := new_message("/address/test")
			msg.append(int32(1122))
			msg.append(stringArgument)
			if err := client.Send(msg); err != nil {
				t.Error(err)
				done.Done()
				done.Done()
				return
			}
		}

		done.Done()

		select {
		case <-timeout:
		case <-finish:
		}
		done.Done()
	}()

	done.Wait()
}

fn server_message_dispatching_udp_test() {
	// Attempting to send a message larger than this (the exact threshold depends
	// on your OS, etc.) results in an error like:
	//
	//   write udp 127.0.0.1:52496->127.0.0.1:6677: write: message too long
	//
	// This is expected for UDP. The practical guaranteed packet size limit for
	// UDP is 576 bytes, and some of that is taken up by protocol overhead.
	//
	// Reference:
	// https://forum.juce.com/t/osc-blobs-are-lost-above-certain-size/20241/2
	testServerMessageDispatching(t, randomString(500))
}

fn server_message_receiving_test(stringArgument string) {
	port := 6677

	finish := make(chan bool)
	start := make(chan bool)
	done := sync.WaitGroup{}
	done.Add(2)

	// Start the server in a go-routine
	go func() {
		server := &Server{}

		c, err := net.ListenPacket("udp", "localhost:"+strconv.Itoa(port))
		if err != nil {
			t.Error(err)
			return
		}
		defer c.Close()

		// Start the client
		start <- true

		packet, err := server.ReceivePacket(c)
		if err != nil {
			t.Errorf("server error: %v", err)
			return
		}
		if packet == nil {
			t.Error("nil packet")
			return
		}

		msg := packet.(*Message)
		if msg.CountArguments() != 3 {
			t.Errorf("Argument length should be 3 and is: %d\n", msg.CountArguments())
		}
		if msg.Arguments[0].(int32) != 1122 {
			t.Error("Argument should be 1122 and is: " + string(msg.Arguments[0].(int32)))
		}
		if msg.Arguments[1].(int32) != 3344 {
			t.Error("Argument should be 3344 and is: " + string(msg.Arguments[1].(int32)))
		}

		receivedString := msg.Arguments[2].(string)
		if len(receivedString) != len(stringArgument) {
			t.Errorf(
				"String argument length should be %d and is %d",
				len(stringArgument),
				len(receivedString),
			)
		} else if receivedString != stringArgument {
			t.Errorf(
				"Argument should be %s and is: %s", stringArgument, receivedString,
			)
		}

		c.Close()
		finish <- true
	}()

	go func() {
		timeout := time.After(5 * time.Second)
		select {
		case <-timeout:
		case <-start:
			client := NewClient("localhost", port)
			msg := new_message("/address/test")
			msg.append(int32(1122))
			msg.append(int32(3344))
			msg.append(stringArgument)
			time.Sleep(500 * time.Millisecond)
			if err := client.Send(msg); err != nil {
				t.Error(err)
				done.Done()
				done.Done()
				return
			}
		}

		done.Done()

		select {
		case <-timeout:
		case <-finish:
		}
		done.Done()
	}()

	done.Wait()
}

// source: https://www.calhoun.io/creating-random-strings-in-go/
fn random_string(length int) string {
	const charset = "abcdefghijklmnopqrstuvwxyzABCDEFGHIJKLMNOPQRSTUVWXYZ"
	var seededRand = rand.New(rand.NewSource(time.Now().UnixNano()))

	b := make([]byte, length)
	for i := range b {
		b[i] = charset[seededRand.Intn(len(charset))]
	}
	return string(b)
}

fn server_message_receiving_udp_test() {
	// Attempting to send a message larger than this (the exact threshold depends
	// on your OS, etc.) results in an error like:
	//
	//   write udp 127.0.0.1:52496->127.0.0.1:6677: write: message too long
	//
	// This is expected for UDP. The practical guaranteed packet size limit for
	// UDP is 576 bytes, and some of that is taken up by protocol overhead.
	//
	// Reference:
	// https://forum.juce.com/t/osc-blobs-are-lost-above-certain-size/20241/2
	testServerMessageReceiving(t, randomString(500))
}

fn read_timeout_test() {
	start := make(chan bool)
	wg := sync.WaitGroup{}
	wg.Add(2)

	go func() {
		defer wg.Done()

		select {
		case <-time.After(5 * time.Second):
			t.Error("timed out")
			wg.Done()
		case <-start:
			client := NewClient("localhost", 6677)
			msg := new_message("/address/test1")
			err := client.Send(msg)
			if err != nil {
				t.Error(err)
			}

			time.Sleep(500 * time.Millisecond)
			msg = new_message("/address/test2")
			err = client.Send(msg)
			if err != nil {
				t.Error(err)
			}
		}
	}()

	go func() {
		defer wg.Done()

		server := &Server{ReadTimeout: 300 * time.Millisecond}
		c, err := net.ListenPacket("udp", "localhost:6677")
		if err != nil {
			t.Error(err)
		}
		defer c.Close()

		// Start the client
		start <- true
		p, err := server.ReceivePacket(c)
		if err != nil {
			t.Errorf("server error: %v", err)
			return
		}
		if got, want := p.(*Message).Address, "/address/test1"; got != want {
			t.Errorf("wrong address; got = %s, want = %s", got, want)
			return
		}

		// Second receive should time out since client is delayed 150 milliseconds
		if _, err = server.ReceivePacket(c); err == nil {
			t.Errorf("expected error")
			return
		}

		// Next receive should get it
		p, err = server.ReceivePacket(c)
		if err != nil {
			t.Errorf("server error: %v", err)
			return
		}
		if got, want := p.(*Message).Address, "/address/test2"; got != want {
			t.Errorf("wrong address; got = %s, want = %s", got, want)
			return
		}
	}()

	wg.Wait()
}

fn read_blob_test() {
	for _, tt := range []struct {
		name    string
		args    []byte
		want    []byte
		want1   int
		wantErr bool
	}{
		{"negative value", []byte{255, 255, 255, 255}, nil, 0, true},
		{"large value", []byte{0, 1, 17, 112}, nil, 0, true},
		{"regular value", []byte{0, 0, 0, 1, 10, 0, 0, 0}, []byte{10}, 8, false},
	} {
		t.Run(tt.name, func() {
			got, got1, err := readBlob(bufio.NewReader(bytes.NewBuffer(tt.args)))
			if (err != nil) != tt.wantErr {
				t.Errorf("readBlob() error = %v, wantErr %v", err, tt.wantErr)
				return
			}
			if !reflect.DeepEqual(got, tt.want) {
				t.Errorf("readBlob() got = %v, want %v", got, tt.want)
			}
			if got1 != tt.want1 {
				t.Errorf("readBlob() got1 = %v, want %v", got1, tt.want1)
			}
		})
	}
}

fn read_padded_string_test() {
	for _, tt := range []struct {
		buf []byte // buffer
		n   int    // bytes needed
		s   string // resulting string
		e   error  // expected error
	}{
		{[]byte{'t', 'e', 's', 't', 'S', 't', 'r', 'i', 'n', 'g', 0, 0}, 12, "testString", nil},
		{[]byte{'t', 'e', 's', 't', 'e', 'r', 's', 0}, 8, "testers", nil},
		{[]byte{'t', 'e', 's', 't', 's', 0, 0, 0}, 8, "tests", nil},
		{[]byte{'t', 'e', 's', 't', 0, 0, 0, 0}, 8, "test", nil},
		{[]byte{}, 0, "", io.EOF},
		{[]byte{'t', 'e', 's', 0}, 4, "tes", nil},             // OSC uses null terminated strings
		{[]byte{'t', 'e', 's', 0, 0, 0, 0, 0}, 4, "tes", nil}, // Additional nulls should be ignored
		{[]byte{'t', 'e', 's', 0, 0, 0}, 4, "tes", nil},       // Whether or not the nulls fall on a 4 byte padding boundary
		{[]byte{'t', 'e', 's', 't'}, 0, "", io.EOF},           // if there is no null byte at the end, it doesn't work.
	} {
		buf := bytes.NewBuffer(tt.buf)
		s, n, err := readPaddedString(bufio.NewReader(buf))
		if got, want := err, tt.e; got != want {
			t.Errorf("%q: Unexpected error reading padded string; got = %q, want = %q", tt.s, got, want)
		}
		if got, want := n, tt.n; got != want {
			t.Errorf("%q: Bytes needed don't match; got = %d, want = %d", tt.s, got, want)
		}
		if got, want := s, tt.s; got != want {
			t.Errorf("%q: Strings don't match; got = %q, want = %q", tt.s, got, want)
		}
	}
}

fn write_padded_string_test() {
	for _, tt := range []struct {
		s   string // string
		buf []byte // resulting buffer
		n   int    // bytes expected
	}{
		{"testString", []byte{'t', 'e', 's', 't', 'S', 't', 'r', 'i', 'n', 'g', 0, 0}, 12},
		{"testers", []byte{'t', 'e', 's', 't', 'e', 'r', 's', 0}, 8},
		{"tests", []byte{'t', 'e', 's', 't', 's', 0, 0, 0}, 8},
		{"test", []byte{'t', 'e', 's', 't', 0, 0, 0, 0}, 8},
		{"tes", []byte{'t', 'e', 's', 0}, 4},
		{"tes\x00", []byte{'t', 'e', 's', 0}, 4},                 // Don't add a second null terminator if one is already present
		{"tes\x00\x00\x00\x00\x00", []byte{'t', 'e', 's', 0}, 4}, // Skip extra nulls
		{"tes\x00\x00\x00", []byte{'t', 'e', 's', 0}, 4},         // Even if they don't fall on a 4 byte padding boundary
		{"", []byte{0, 0, 0, 0}, 4},                              // OSC uses null terminated strings, padded to the 4 byte boundary
	} {
		buf := []byte{}
		bytesBuffer := bytes.NewBuffer(buf)

		n, err := writePaddedString(tt.s, bytesBuffer)
		if err != nil {
			t.Errorf(err.Error())
		}
		if got, want := n, tt.n; got != want {
			t.Errorf("%q: Count of bytes written don't match; got = %d, want = %d", tt.s, got, want)
		}
		if got, want := bytesBuffer, tt.buf; !bytes.Equal(got.Bytes(), want) {
			t.Errorf("%q: Buffers don't match; got = %q, want = %q", tt.s, got.Bytes(), want)
		}
	}
}

fn pad_bytes_needed_test() {
	var n int
	n = padBytesNeeded(4)
	if n != 0 {
		t.Errorf("Number of pad bytes should be 0 and is: %d", n)
	}

	n = padBytesNeeded(3)
	if n != 1 {
		t.Errorf("Number of pad bytes should be 1 and is: %d", n)
	}

	n = padBytesNeeded(2)
	if n != 2 {
		t.Errorf("Number of pad bytes should be 2 and is: %d", n)
	}

	n = padBytesNeeded(1)
	if n != 3 {
		t.Errorf("Number of pad bytes should be 3 and is: %d", n)
	}

	n = padBytesNeeded(0)
	if n != 0 {
		t.Errorf("Number of pad bytes should be 0 and is: %d", n)
	}

	n = padBytesNeeded(5)
	if n != 3 {
		t.Errorf("Number of pad bytes should be 3 and is: %d", n)
	}

	n = padBytesNeeded(7)
	if n != 1 {
		t.Errorf("Number of pad bytes should be 1 and is: %d", n)
	}

	n = padBytesNeeded(32)
	if n != 0 {
		t.Errorf("Number of pad bytes should be 0 and is: %d", n)
	}

	n = padBytesNeeded(63)
	if n != 1 {
		t.Errorf("Number of pad bytes should be 1 and is: %d", n)
	}

	n = padBytesNeeded(10)
	if n != 2 {
		t.Errorf("Number of pad bytes should be 2 and is: %d", n)
	}
}

fn type_tags_string_test() {
	msg := new_message("/some/address")
	msg.append(int32(100))
	msg.append(true)
	msg.append(false)

	typeTags, err := msg.TypeTags()
	if err != nil {
		t.Error(err.Error())
	}

	if typeTags != ",iTF" {
		t.Errorf("Type tag string should be ',iTF' and is: %s", typeTags)
	}
}

fn client_set_local_addr_test() {
	client := NewClient("localhost", 8967)
	err := client.SetLocalAddr("localhost", 41789)
	if err != nil {
		t.Error(err.Error())
	}
	expectedAddr := "127.0.0.1:41789"
	if client.laddr.String() != expectedAddr {
		t.Errorf("Expected laddr to be %s but was %s", expectedAddr, client.laddr.String())
	}
}

fn parse_packet_test() {
	for _, tt := range []struct {
		desc string
		msg  string
		pkt  Packet
		ok   bool
	}{
		{"no_args",
			"/a/b/c" + nulls(2) + "," + nulls(3),
			makePacket("/a/b/c", nil),
			true},
		{"string_arg",
			"/d/e/f" + nulls(2) + ",s" + nulls(2) + "foo" + nulls(1),
			makePacket("/d/e/f", []string{"foo"}),
			true},
		{"empty", "", nil, false},
	} {
		pkt, err := ParsePacket(tt.msg)
		if err != nil && tt.ok {
			t.Errorf("%s: ParsePacket() returned unexpected error; %s", tt.desc, err)
		}
		if err == nil && !tt.ok {
			t.Errorf("%s: ParsePacket() expected error", tt.desc)
		}
		if !tt.ok {
			continue
		}

		pktBytes, err := pkt.MarshalBinary()
		if err != nil {
			t.Errorf("%s: failure converting pkt to byte array; %s", tt.desc, err)
			continue
		}
		ttpktBytes, err := tt.pkt.MarshalBinary()
		if err != nil {
			t.Errorf("%s: failure converting tt.pkt to byte array; %s", tt.desc, err)
			continue
		}
		if got, want := pktBytes, ttpktBytes; !reflect.DeepEqual(got, want) {
			t.Errorf("%s: ParsePacket() as bytes = '%s', want = '%s'", tt.desc, got, want)
			continue
		}
	}
}

fn osc_message_match_test() {
	tc := []struct {
		desc        string
		addr        string
		addrPattern string
		want        bool
	}{
		{
			"match everything",
			"*",
			"/a/b",
			true,
		},
		{
			"don't match",
			"/a/b",
			"/a",
			false,
		},
		{
			"match alternatives",
			"/a/{foo,bar}",
			"/a/foo",
			true,
		},
		{
			"don't match if address is not part of the alternatives",
			"/a/{foo,bar}",
			"/a/bob",
			false,
		},
	}

	for _, tt := range tc {
		msg := new_message(tt.addr)

		got := msg.Match(tt.addrPattern)
		if got != tt.want {
			t.Errorf("%s: msg.Match('%s') = '%t', want = '%t'", tt.desc, tt.addrPattern, got, tt.want)
		}
	}
}

fn time_to_timetag_test() {
	tc := []struct {
		desc  string
		input time.Time
		want  uint64
	}{
		{
			"return zero time instance when timetag = 1",
			time.Time{},
			1,
		},
		{
			"calculate correct timetag without parts of second",
			time.Unix(1646694561, 0),
			16560033939226361856,
		},
		{
			"calculate correct timetag with parts of second",
			time.Unix(1646694561, 500),
			16560033939226364003,
		},
	}

	for _, tt := range tc {
		got := timeToTimetag(tt.input)
		if got != tt.want {
			t.Errorf("%s: timeToTimetag: '%d', want = '%d'", tt.desc, got, tt.want)
		}
	}
}

fn timetag_to_time_test() {
	tc := []struct {
		desc  string
		input uint64
		want  time.Time
	}{
		{
			"return zero time instance when timetag = 1",
			1,
			time.Time{},
		},
		{
			"calculate correct timetag without parts of second",
			16560033939226361856,
			time.Unix(1646694561, 0),
		},
		{
			"calculate correct timetag with parts of second",
			16560033939226364004,
			time.Unix(1646694561, 500),
		},
	}

	for _, tt := range tc {
		got := timetagToTime(tt.input)
		if got != tt.want {
			t.Errorf("%s: timetagToTime: '%v', want = '%v'", tt.desc, got, tt.want)
		}
	}
}

const zero = string(byte(0))

// nulls returns a string of `i` nulls.
fn nulls(i int) string {
	s := ""
	for j := 0; j < i; j++ {
		s += zero
	}
	return s
}

// makePacket creates a fake Message Packet.
fn make_packet(addr string, args []string) Packet {
	msg := new_message(addr)
	for _, arg := range args {
		msg.append(arg)
	}
	return msg
}
